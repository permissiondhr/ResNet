module bn_res
#(
    parameter DATA_WIDTH   = 16,
    parameter PARA_WIDTH   = 16,
    parameter CHANNEL_NUM  = 128,
	parameter FM_DEPTH	   = 64
)
(
    // GLOBAL SIGNALS
    input   wire                    			clk             ,    			// System Clock
    input   wire                    			rstn            ,    			// System Reset, Active LOW
    input   wire                    			data_in_valid   ,    			// DATA Enable signal, Active HIGH
    input   wire signed [PARA_WIDTH - 1 : 0] 	bn_a     [CHANNEL_NUM - 1 : 0],	// Parameter of BN
    input   wire signed [PARA_WIDTH - 1 : 0] 	bn_b     [CHANNEL_NUM - 1 : 0],	// Parameter of BN
    input   wire signed [DATA_WIDTH - 1 : 0] 	res      [FM_DEPTH - 1    : 0],	// Residual
    input   wire signed [5 : 0] 				data_in  [CHANNEL_NUM - 1 : 0],	// Data from partial_sum
    output  wire signed [DATA_WIDTH - 1 : 0] 	data_out [CHANNEL_NUM - 1 : 0],	// Data to RPReLU
    output  reg                     			data_out_valid              	// DATA Enable signal to RPReLU
);

reg  signed [PARA_WIDTH + DATA_WIDTH -1: 0] product [CHANNEL_NUM - 1 : 0];
wire signed [DATA_WIDTH - 1 : 0] 			data_in_extended [CHANNEL_NUM - 1 : 0];
wire signed [PARA_WIDTH + DATA_WIDTH -1: 0]	product_sr [CHANNEL_NUM - 1 : 0];

genvar i;
generate
	for(i = 0; i < CHANNEL_NUM; i = i + 1) begin
		assign data_in_extended[i] = {{10{data_in[i][5]}}, data_in[i]};
		always @(posedge clk or negedge rstn) begin    
	        if(~rstn) begin
	            data_out_valid  <= 0;
	            product[i] 		<= 0;
	        end 
			else begin
				if(data_in_valid) begin
	            	data_out_valid  <= 1;
	            	product[i] 		<= bn_a[i] * data_in_extended[i];
	        	end 
				else begin
	            	data_out_valid  <= 0;
	            	product[i] 		<= product[i];
				end
	        end
	    end

		assign product_sr[i] = product[i] >>> 8;

		if (i < FM_DEPTH)
			assign data_out[i] = product_sr[i] + bn_b[i]  + res[i];
		else
			assign data_out[i] = product_sr[i] + bn_b[i];
	end
endgenerate

endmodule // bn_res_layer4